* Inductances
L0	2	9
L1	2	14
L2	9	7
L3	9	4
L4	14	16
L5	7	3
L6	7	10
L7	4	3
L8	4	6
L9	3	13

* Ports
P1+ NbN2	16	0
P2+ NbN2	10	0
P3+ NbN2	13	0
P4+ NbN2	6	0
.end